
my first comment
my second comment
